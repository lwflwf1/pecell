/home/wyc/Project/To_Vrf/rtl/pe_rram.sv